module cos_generator (
    input  wire [7:0] address,  // ??a ch? 8-bit
    input  wire       clock,    // Clock
    output reg  [7:0] q         // Gi� tr? COS ??u ra
);

reg [7:0] cos_lut [0:255]; // Look-Up Table 256 gi� tr?

initial begin
    // Kh?i t?o LUT v?i gi� tr? COS (gi? s? bi�n ?? 127, offset 128)
cos_lut[0] = 8'd255;
cos_lut[1] = 8'd255;
cos_lut[2] = 8'd255;
cos_lut[3] = 8'd255;
cos_lut[4] = 8'd254;
cos_lut[5] = 8'd254;
cos_lut[6] = 8'd254;
cos_lut[7] = 8'd253;
cos_lut[8] = 8'd253;
cos_lut[9] = 8'd252;
cos_lut[10] = 8'd251;
cos_lut[11] = 8'd250;
cos_lut[12] = 8'd250;
cos_lut[13] = 8'd249;
cos_lut[14] = 8'd248;
cos_lut[15] = 8'd246;
cos_lut[16] = 8'd245;
cos_lut[17] = 8'd244;
cos_lut[18] = 8'd243;
cos_lut[19] = 8'd241;
cos_lut[20] = 8'd240;
cos_lut[21] = 8'd239;
cos_lut[22] = 8'd237;
cos_lut[23] = 8'd235;
cos_lut[24] = 8'd234;
cos_lut[25] = 8'd232;
cos_lut[26] = 8'd230;
cos_lut[27] = 8'd228;
cos_lut[28] = 8'd226;
cos_lut[29] = 8'd224;
cos_lut[30] = 8'd222;
cos_lut[31] = 8'd220;
cos_lut[32] = 8'd218;
cos_lut[33] = 8'd216;
cos_lut[34] = 8'd213;
cos_lut[35] = 8'd211;
cos_lut[36] = 8'd209;
cos_lut[37] = 8'd206;
cos_lut[38] = 8'd204;
cos_lut[39] = 8'd201;
cos_lut[40] = 8'd199;
cos_lut[41] = 8'd196;
cos_lut[42] = 8'd193;
cos_lut[43] = 8'd191;
cos_lut[44] = 8'd188;
cos_lut[45] = 8'd185;
cos_lut[46] = 8'd182;
cos_lut[47] = 8'd179;
cos_lut[48] = 8'd177;
cos_lut[49] = 8'd174;
cos_lut[50] = 8'd171;
cos_lut[51] = 8'd168;
cos_lut[52] = 8'd165;
cos_lut[53] = 8'd162;
cos_lut[54] = 8'd159;
cos_lut[55] = 8'd156;
cos_lut[56] = 8'd153;
cos_lut[57] = 8'd150;
cos_lut[58] = 8'd147;
cos_lut[59] = 8'd144;
cos_lut[60] = 8'd140;
cos_lut[61] = 8'd137;
cos_lut[62] = 8'd134;
cos_lut[63] = 8'd131;
cos_lut[64] = 8'd128;
cos_lut[65] = 8'd125;
cos_lut[66] = 8'd122;
cos_lut[67] = 8'd119;
cos_lut[68] = 8'd116;
cos_lut[69] = 8'd112;
cos_lut[70] = 8'd109;
cos_lut[71] = 8'd106;
cos_lut[72] = 8'd103;
cos_lut[73] = 8'd100;
cos_lut[74] = 8'd97;
cos_lut[75] = 8'd94;
cos_lut[76] = 8'd91;
cos_lut[77] = 8'd88;
cos_lut[78] = 8'd85;
cos_lut[79] = 8'd82;
cos_lut[80] = 8'd79;
cos_lut[81] = 8'd77;
cos_lut[82] = 8'd74;
cos_lut[83] = 8'd71;
cos_lut[84] = 8'd68;
cos_lut[85] = 8'd65;
cos_lut[86] = 8'd63;
cos_lut[87] = 8'd60;
cos_lut[88] = 8'd57;
cos_lut[89] = 8'd55;
cos_lut[90] = 8'd52;
cos_lut[91] = 8'd50;
cos_lut[92] = 8'd47;
cos_lut[93] = 8'd45;
cos_lut[94] = 8'd43;
cos_lut[95] = 8'd40;
cos_lut[96] = 8'd38;
cos_lut[97] = 8'd36;
cos_lut[98] = 8'd34;
cos_lut[99] = 8'd32;
cos_lut[100] = 8'd30;
cos_lut[101] = 8'd28;
cos_lut[102] = 8'd26;
cos_lut[103] = 8'd24;
cos_lut[104] = 8'd22;
cos_lut[105] = 8'd21;
cos_lut[106] = 8'd19;
cos_lut[107] = 8'd17;
cos_lut[108] = 8'd16;
cos_lut[109] = 8'd15;
cos_lut[110] = 8'd13;
cos_lut[111] = 8'd12;
cos_lut[112] = 8'd11;
cos_lut[113] = 8'd10;
cos_lut[114] = 8'd8;
cos_lut[115] = 8'd7;
cos_lut[116] = 8'd6;
cos_lut[117] = 8'd6;
cos_lut[118] = 8'd5;
cos_lut[119] = 8'd4;
cos_lut[120] = 8'd3;
cos_lut[121] = 8'd3;
cos_lut[122] = 8'd2;
cos_lut[123] = 8'd2;
cos_lut[124] = 8'd2;
cos_lut[125] = 8'd1;
cos_lut[126] = 8'd1;
cos_lut[127] = 8'd1;
cos_lut[128] = 8'd1;
cos_lut[129] = 8'd1;
cos_lut[130] = 8'd1;
cos_lut[131] = 8'd1;
cos_lut[132] = 8'd2;
cos_lut[133] = 8'd2;
cos_lut[134] = 8'd2;
cos_lut[135] = 8'd3;
cos_lut[136] = 8'd3;
cos_lut[137] = 8'd4;
cos_lut[138] = 8'd5;
cos_lut[139] = 8'd6;
cos_lut[140] = 8'd6;
cos_lut[141] = 8'd7;
cos_lut[142] = 8'd8;
cos_lut[143] = 8'd10;
cos_lut[144] = 8'd11;
cos_lut[145] = 8'd12;
cos_lut[146] = 8'd13;
cos_lut[147] = 8'd15;
cos_lut[148] = 8'd16;
cos_lut[149] = 8'd17;
cos_lut[150] = 8'd19;
cos_lut[151] = 8'd21;
cos_lut[152] = 8'd22;
cos_lut[153] = 8'd24;
cos_lut[154] = 8'd26;
cos_lut[155] = 8'd28;
cos_lut[156] = 8'd30;
cos_lut[157] = 8'd32;
cos_lut[158] = 8'd34;
cos_lut[159] = 8'd36;
cos_lut[160] = 8'd38;
cos_lut[161] = 8'd40;
cos_lut[162] = 8'd43;
cos_lut[163] = 8'd45;
cos_lut[164] = 8'd47;
cos_lut[165] = 8'd50;
cos_lut[166] = 8'd52;
cos_lut[167] = 8'd55;
cos_lut[168] = 8'd57;
cos_lut[169] = 8'd60;
cos_lut[170] = 8'd63;
cos_lut[171] = 8'd65;
cos_lut[172] = 8'd68;
cos_lut[173] = 8'd71;
cos_lut[174] = 8'd74;
cos_lut[175] = 8'd77;
cos_lut[176] = 8'd79;
cos_lut[177] = 8'd82;
cos_lut[178] = 8'd85;
cos_lut[179] = 8'd88;
cos_lut[180] = 8'd91;
cos_lut[181] = 8'd94;
cos_lut[182] = 8'd97;
cos_lut[183] = 8'd100;
cos_lut[184] = 8'd103;
cos_lut[185] = 8'd106;
cos_lut[186] = 8'd109;
cos_lut[187] = 8'd112;
cos_lut[188] = 8'd116;
cos_lut[189] = 8'd119;
cos_lut[190] = 8'd122;
cos_lut[191] = 8'd125;
cos_lut[192] = 8'd128;
cos_lut[193] = 8'd131;
cos_lut[194] = 8'd134;
cos_lut[195] = 8'd137;
cos_lut[196] = 8'd140;
cos_lut[197] = 8'd144;
cos_lut[198] = 8'd147;
cos_lut[199] = 8'd150;
cos_lut[200] = 8'd153;
cos_lut[201] = 8'd156;
cos_lut[202] = 8'd159;
cos_lut[203] = 8'd162;
cos_lut[204] = 8'd165;
cos_lut[205] = 8'd168;
cos_lut[206] = 8'd171;
cos_lut[207] = 8'd174;
cos_lut[208] = 8'd177;
cos_lut[209] = 8'd179;
cos_lut[210] = 8'd182;
cos_lut[211] = 8'd185;
cos_lut[212] = 8'd188;
cos_lut[213] = 8'd191;
cos_lut[214] = 8'd193;
cos_lut[215] = 8'd196;
cos_lut[216] = 8'd199;
cos_lut[217] = 8'd201;
cos_lut[218] = 8'd204;
cos_lut[219] = 8'd206;
cos_lut[220] = 8'd209;
cos_lut[221] = 8'd211;
cos_lut[222] = 8'd213;
cos_lut[223] = 8'd216;
cos_lut[224] = 8'd218;
cos_lut[225] = 8'd220;
cos_lut[226] = 8'd222;
cos_lut[227] = 8'd224;
cos_lut[228] = 8'd226;
cos_lut[229] = 8'd228;
cos_lut[230] = 8'd230;
cos_lut[231] = 8'd232;
cos_lut[232] = 8'd234;
cos_lut[233] = 8'd235;
cos_lut[234] = 8'd237;
cos_lut[235] = 8'd239;
cos_lut[236] = 8'd240;
cos_lut[237] = 8'd241;
cos_lut[238] = 8'd243;
cos_lut[239] = 8'd244;
cos_lut[240] = 8'd245;
cos_lut[241] = 8'd246;
cos_lut[242] = 8'd248;
cos_lut[243] = 8'd249;
cos_lut[244] = 8'd250;
cos_lut[245] = 8'd250;
cos_lut[246] = 8'd251;
cos_lut[247] = 8'd252;
cos_lut[248] = 8'd253;
cos_lut[249] = 8'd253;
cos_lut[250] = 8'd254;
cos_lut[251] = 8'd254;
cos_lut[252] = 8'd254;
cos_lut[253] = 8'd255;
cos_lut[254] = 8'd255;
cos_lut[255] = 8'd255;
end

always @(posedge clock) begin
    q <= cos_lut[address]; // L?y gi� tr? t? LUT theo ??a ch?
end

endmodule
