module sin_generator (
    input  wire [7:0] address,  
    input  wire       clock,    
    output reg  [7:0] q        
);

reg [7:0] sin_lut [0:255]; 

initial begin
sin_lut[0] = 8'h00;
sin_lut[1] = 8'h01;
sin_lut[2] = 8'h02;
sin_lut[3] = 8'h03;
sin_lut[4] = 8'h04;
sin_lut[5] = 8'h05;
sin_lut[6] = 8'h06;
sin_lut[7] = 8'h07;
sin_lut[8] = 8'h08;
sin_lut[9] = 8'h09;
sin_lut[10] = 8'h0A;
sin_lut[11] = 8'h0B;
sin_lut[12] = 8'h0C;
sin_lut[13] = 8'h0D;
sin_lut[14] = 8'h0E;
sin_lut[15] = 8'h0F;
sin_lut[16] = 8'h10;
sin_lut[17] = 8'h11;
sin_lut[18] = 8'h12;
sin_lut[19] = 8'h13;
sin_lut[20] = 8'h14;
sin_lut[21] = 8'h15;
sin_lut[22] = 8'h16;
sin_lut[23] = 8'h16;
sin_lut[24] = 8'h17;
sin_lut[25] = 8'h18;
sin_lut[26] = 8'h19;
sin_lut[27] = 8'h1A;
sin_lut[28] = 8'h1B;
sin_lut[29] = 8'h1B;
sin_lut[30] = 8'h1C;
sin_lut[31] = 8'h1D;
sin_lut[32] = 8'h1E;
sin_lut[33] = 8'h1E;
sin_lut[34] = 8'h1F;
sin_lut[35] = 8'h20;
sin_lut[36] = 8'h20;
sin_lut[37] = 8'h21;
sin_lut[38] = 8'h22;
sin_lut[39] = 8'h22;
sin_lut[40] = 8'h23;
sin_lut[41] = 8'h23;
sin_lut[42] = 8'h24;
sin_lut[43] = 8'h25;
sin_lut[44] = 8'h25;
sin_lut[45] = 8'h26;
sin_lut[46] = 8'h26;
sin_lut[47] = 8'h26;
sin_lut[48] = 8'h27;
sin_lut[49] = 8'h27;
sin_lut[50] = 8'h28;
sin_lut[51] = 8'h28;
sin_lut[52] = 8'h28;
sin_lut[53] = 8'h28;
sin_lut[54] = 8'h29;
sin_lut[55] = 8'h29;
sin_lut[56] = 8'h29;
sin_lut[57] = 8'h29;
sin_lut[58] = 8'h2A;
sin_lut[59] = 8'h2A;
sin_lut[60] = 8'h2A;
sin_lut[61] = 8'h2A;
sin_lut[62] = 8'h2A;
sin_lut[63] = 8'h2A;
sin_lut[64] = 8'h2A;
sin_lut[65] = 8'h2A;
sin_lut[66] = 8'h2A;
sin_lut[67] = 8'h2A;
sin_lut[68] = 8'h2A;
sin_lut[69] = 8'h2A;
sin_lut[70] = 8'h2A;
sin_lut[71] = 8'h29;
sin_lut[72] = 8'h29;
sin_lut[73] = 8'h29;
sin_lut[74] = 8'h29;
sin_lut[75] = 8'h28;
sin_lut[76] = 8'h28;
sin_lut[77] = 8'h28;
sin_lut[78] = 8'h28;
sin_lut[79] = 8'h27;
sin_lut[80] = 8'h27;
sin_lut[81] = 8'h26;
sin_lut[82] = 8'h26;
sin_lut[83] = 8'h26;
sin_lut[84] = 8'h25;
sin_lut[85] = 8'h25;
sin_lut[86] = 8'h24;
sin_lut[87] = 8'h23;
sin_lut[88] = 8'h23;
sin_lut[89] = 8'h22;
sin_lut[90] = 8'h22;
sin_lut[91] = 8'h21;
sin_lut[92] = 8'h20;
sin_lut[93] = 8'h20;
sin_lut[94] = 8'h1F;
sin_lut[95] = 8'h1E;
sin_lut[96] = 8'h1E;
sin_lut[97] = 8'h1D;
sin_lut[98] = 8'h1C;
sin_lut[99] = 8'h1B;
sin_lut[100] = 8'h1B;
sin_lut[101] = 8'h1A;
sin_lut[102] = 8'h19;
sin_lut[103] = 8'h18;
sin_lut[104] = 8'h17;
sin_lut[105] = 8'h16;
sin_lut[106] = 8'h16;
sin_lut[107] = 8'h15;
sin_lut[108] = 8'h14;
sin_lut[109] = 8'h13;
sin_lut[110] = 8'h12;
sin_lut[111] = 8'h11;
sin_lut[112] = 8'h10;
sin_lut[113] = 8'h0F;
sin_lut[114] = 8'h0E;
sin_lut[115] = 8'h0D;
sin_lut[116] = 8'h0C;
sin_lut[117] = 8'h0B;
sin_lut[118] = 8'h0A;
sin_lut[119] = 8'h09;
sin_lut[120] = 8'h08;
sin_lut[121] = 8'h07;
sin_lut[122] = 8'h06;
sin_lut[123] = 8'h05;
sin_lut[124] = 8'h04;
sin_lut[125] = 8'h03;
sin_lut[126] = 8'h02;
sin_lut[127] = 8'h01;
sin_lut[128] = 8'h00;
sin_lut[129] = 8'hFF;
sin_lut[130] = 8'hFE;
sin_lut[131] = 8'hFD;
sin_lut[132] = 8'hFC;
sin_lut[133] = 8'hFB;
sin_lut[134] = 8'hFA;
sin_lut[135] = 8'hF9;
sin_lut[136] = 8'hF8;
sin_lut[137] = 8'hF7;
sin_lut[138] = 8'hF6;
sin_lut[139] = 8'hF5;
sin_lut[140] = 8'hF4;
sin_lut[141] = 8'hF3;
sin_lut[142] = 8'hF2;
sin_lut[143] = 8'hF1;
sin_lut[144] = 8'hF0;
sin_lut[145] = 8'hEF;
sin_lut[146] = 8'hEE;
sin_lut[147] = 8'hED;
sin_lut[148] = 8'hEC;
sin_lut[149] = 8'hEB;
sin_lut[150] = 8'hEA;
sin_lut[151] = 8'hEA;
sin_lut[152] = 8'hE9;
sin_lut[153] = 8'hE8;
sin_lut[154] = 8'hE7;
sin_lut[155] = 8'hE6;
sin_lut[156] = 8'hE5;
sin_lut[157] = 8'hE5;
sin_lut[158] = 8'hE4;
sin_lut[159] = 8'hE3;
sin_lut[160] = 8'hE2;
sin_lut[161] = 8'hE2;
sin_lut[162] = 8'hE1;
sin_lut[163] = 8'hE0;
sin_lut[164] = 8'hE0;
sin_lut[165] = 8'hDF;
sin_lut[166] = 8'hDE;
sin_lut[167] = 8'hDE;
sin_lut[168] = 8'hDD;
sin_lut[169] = 8'hDD;
sin_lut[170] = 8'hDC;
sin_lut[171] = 8'hDB;
sin_lut[172] = 8'hDB;
sin_lut[173] = 8'hDA;
sin_lut[174] = 8'hDA;
sin_lut[175] = 8'hDA;
sin_lut[176] = 8'hD9;
sin_lut[177] = 8'hD9;
sin_lut[178] = 8'hD8;
sin_lut[179] = 8'hD8;
sin_lut[180] = 8'hD8;
sin_lut[181] = 8'hD8;
sin_lut[182] = 8'hD7;
sin_lut[183] = 8'hD7;
sin_lut[184] = 8'hD7;
sin_lut[185] = 8'hD7;
sin_lut[186] = 8'hD6;
sin_lut[187] = 8'hD6;
sin_lut[188] = 8'hD6;
sin_lut[189] = 8'hD6;
sin_lut[190] = 8'hD6;
sin_lut[191] = 8'hD6;
sin_lut[192] = 8'hD6;
sin_lut[193] = 8'hD6;
sin_lut[194] = 8'hD6;
sin_lut[195] = 8'hD6;
sin_lut[196] = 8'hD6;
sin_lut[197] = 8'hD6;
sin_lut[198] = 8'hD6;
sin_lut[199] = 8'hD7;
sin_lut[200] = 8'hD7;
sin_lut[201] = 8'hD7;
sin_lut[202] = 8'hD7;
sin_lut[203] = 8'hD8;
sin_lut[204] = 8'hD8;
sin_lut[205] = 8'hD8;
sin_lut[206] = 8'hD8;
sin_lut[207] = 8'hD9;
sin_lut[208] = 8'hD9;
sin_lut[209] = 8'hDA;
sin_lut[210] = 8'hDA;
sin_lut[211] = 8'hDA;
sin_lut[212] = 8'hDB;
sin_lut[213] = 8'hDB;
sin_lut[214] = 8'hDC;
sin_lut[215] = 8'hDD;
sin_lut[216] = 8'hDD;
sin_lut[217] = 8'hDE;
sin_lut[218] = 8'hDE;
sin_lut[219] = 8'hDF;
sin_lut[220] = 8'hE0;
sin_lut[221] = 8'hE0;
sin_lut[222] = 8'hE1;
sin_lut[223] = 8'hE2;
sin_lut[224] = 8'hE2;
sin_lut[225] = 8'hE3;
sin_lut[226] = 8'hE4;
sin_lut[227] = 8'hE5;
sin_lut[228] = 8'hE5;
sin_lut[229] = 8'hE6;
sin_lut[230] = 8'hE7;
sin_lut[231] = 8'hE8;
sin_lut[232] = 8'hE9;
sin_lut[233] = 8'hEA;
sin_lut[234] = 8'hEA;
sin_lut[235] = 8'hEB;
sin_lut[236] = 8'hEC;
sin_lut[237] = 8'hED;
sin_lut[238] = 8'hEE;
sin_lut[239] = 8'hEF;
sin_lut[240] = 8'hF0;
sin_lut[241] = 8'hF1;
sin_lut[242] = 8'hF2;
sin_lut[243] = 8'hF3;
sin_lut[244] = 8'hF4;
sin_lut[245] = 8'hF5;
sin_lut[246] = 8'hF6;
sin_lut[247] = 8'hF7;
sin_lut[248] = 8'hF8;
sin_lut[249] = 8'hF9;
sin_lut[250] = 8'hFA;
sin_lut[251] = 8'hFB;
sin_lut[252] = 8'hFC;
sin_lut[253] = 8'hFD;
sin_lut[254] = 8'hFE;
sin_lut[255] = 8'hFF;

end

always @(posedge clock) begin
    q <= sin_lut[address]; 
end

endmodule
