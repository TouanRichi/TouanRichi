module cos_generator (
    input  wire [7:0] address,  
    input  wire       clock,    
    output reg  [7:0] q         
);

reg [7:0] cos_lut [0:255]; 

initial begin
cos_lut[0] = 8'h2A;
cos_lut[1] = 8'h2A;
cos_lut[2] = 8'h2A;
cos_lut[3] = 8'h2A;
cos_lut[4] = 8'h2A;
cos_lut[5] = 8'h2A;
cos_lut[6] = 8'h2A;
cos_lut[7] = 8'h29;
cos_lut[8] = 8'h29;
cos_lut[9] = 8'h29;
cos_lut[10] = 8'h29;
cos_lut[11] = 8'h28;
cos_lut[12] = 8'h28;
cos_lut[13] = 8'h28;
cos_lut[14] = 8'h28;
cos_lut[15] = 8'h27;
cos_lut[16] = 8'h27;
cos_lut[17] = 8'h26;
cos_lut[18] = 8'h26;
cos_lut[19] = 8'h26;
cos_lut[20] = 8'h25;
cos_lut[21] = 8'h25;
cos_lut[22] = 8'h24;
cos_lut[23] = 8'h23;
cos_lut[24] = 8'h23;
cos_lut[25] = 8'h22;
cos_lut[26] = 8'h22;
cos_lut[27] = 8'h21;
cos_lut[28] = 8'h20;
cos_lut[29] = 8'h20;
cos_lut[30] = 8'h1F;
cos_lut[31] = 8'h1E;
cos_lut[32] = 8'h1E;
cos_lut[33] = 8'h1D;
cos_lut[34] = 8'h1C;
cos_lut[35] = 8'h1B;
cos_lut[36] = 8'h1B;
cos_lut[37] = 8'h1A;
cos_lut[38] = 8'h19;
cos_lut[39] = 8'h18;
cos_lut[40] = 8'h17;
cos_lut[41] = 8'h16;
cos_lut[42] = 8'h16;
cos_lut[43] = 8'h15;
cos_lut[44] = 8'h14;
cos_lut[45] = 8'h13;
cos_lut[46] = 8'h12;
cos_lut[47] = 8'h11;
cos_lut[48] = 8'h10;
cos_lut[49] = 8'h0F;
cos_lut[50] = 8'h0E;
cos_lut[51] = 8'h0D;
cos_lut[52] = 8'h0C;
cos_lut[53] = 8'h0B;
cos_lut[54] = 8'h0A;
cos_lut[55] = 8'h09;
cos_lut[56] = 8'h08;
cos_lut[57] = 8'h07;
cos_lut[58] = 8'h06;
cos_lut[59] = 8'h05;
cos_lut[60] = 8'h04;
cos_lut[61] = 8'h03;
cos_lut[62] = 8'h02;
cos_lut[63] = 8'h01;
cos_lut[64] = 8'h00;
cos_lut[65] = 8'hFF;
cos_lut[66] = 8'hFE;
cos_lut[67] = 8'hFD;
cos_lut[68] = 8'hFC;
cos_lut[69] = 8'hFB;
cos_lut[70] = 8'hFA;
cos_lut[71] = 8'hF9;
cos_lut[72] = 8'hF8;
cos_lut[73] = 8'hF7;
cos_lut[74] = 8'hF6;
cos_lut[75] = 8'hF5;
cos_lut[76] = 8'hF4;
cos_lut[77] = 8'hF3;
cos_lut[78] = 8'hF2;
cos_lut[79] = 8'hF1;
cos_lut[80] = 8'hF0;
cos_lut[81] = 8'hEF;
cos_lut[82] = 8'hEE;
cos_lut[83] = 8'hED;
cos_lut[84] = 8'hEC;
cos_lut[85] = 8'hEB;
cos_lut[86] = 8'hEA;
cos_lut[87] = 8'hEA;
cos_lut[88] = 8'hE9;
cos_lut[89] = 8'hE8;
cos_lut[90] = 8'hE7;
cos_lut[91] = 8'hE6;
cos_lut[92] = 8'hE5;
cos_lut[93] = 8'hE5;
cos_lut[94] = 8'hE4;
cos_lut[95] = 8'hE3;
cos_lut[96] = 8'hE2;
cos_lut[97] = 8'hE2;
cos_lut[98] = 8'hE1;
cos_lut[99] = 8'hE0;
cos_lut[100] = 8'hE0;
cos_lut[101] = 8'hDF;
cos_lut[102] = 8'hDE;
cos_lut[103] = 8'hDE;
cos_lut[104] = 8'hDD;
cos_lut[105] = 8'hDD;
cos_lut[106] = 8'hDC;
cos_lut[107] = 8'hDB;
cos_lut[108] = 8'hDB;
cos_lut[109] = 8'hDA;
cos_lut[110] = 8'hDA;
cos_lut[111] = 8'hDA;
cos_lut[112] = 8'hD9;
cos_lut[113] = 8'hD9;
cos_lut[114] = 8'hD8;
cos_lut[115] = 8'hD8;
cos_lut[116] = 8'hD8;
cos_lut[117] = 8'hD8;
cos_lut[118] = 8'hD7;
cos_lut[119] = 8'hD7;
cos_lut[120] = 8'hD7;
cos_lut[121] = 8'hD7;
cos_lut[122] = 8'hD6;
cos_lut[123] = 8'hD6;
cos_lut[124] = 8'hD6;
cos_lut[125] = 8'hD6;
cos_lut[126] = 8'hD6;
cos_lut[127] = 8'hD6;
cos_lut[128] = 8'hD6;
cos_lut[129] = 8'hD6;
cos_lut[130] = 8'hD6;
cos_lut[131] = 8'hD6;
cos_lut[132] = 8'hD6;
cos_lut[133] = 8'hD6;
cos_lut[134] = 8'hD6;
cos_lut[135] = 8'hD7;
cos_lut[136] = 8'hD7;
cos_lut[137] = 8'hD7;
cos_lut[138] = 8'hD7;
cos_lut[139] = 8'hD8;
cos_lut[140] = 8'hD8;
cos_lut[141] = 8'hD8;
cos_lut[142] = 8'hD8;
cos_lut[143] = 8'hD9;
cos_lut[144] = 8'hD9;
cos_lut[145] = 8'hDA;
cos_lut[146] = 8'hDA;
cos_lut[147] = 8'hDA;
cos_lut[148] = 8'hDB;
cos_lut[149] = 8'hDB;
cos_lut[150] = 8'hDC;
cos_lut[151] = 8'hDD;
cos_lut[152] = 8'hDD;
cos_lut[153] = 8'hDE;
cos_lut[154] = 8'hDE;
cos_lut[155] = 8'hDF;
cos_lut[156] = 8'hE0;
cos_lut[157] = 8'hE0;
cos_lut[158] = 8'hE1;
cos_lut[159] = 8'hE2;
cos_lut[160] = 8'hE2;
cos_lut[161] = 8'hE3;
cos_lut[162] = 8'hE4;
cos_lut[163] = 8'hE5;
cos_lut[164] = 8'hE5;
cos_lut[165] = 8'hE6;
cos_lut[166] = 8'hE7;
cos_lut[167] = 8'hE8;
cos_lut[168] = 8'hE9;
cos_lut[169] = 8'hEA;
cos_lut[170] = 8'hEA;
cos_lut[171] = 8'hEB;
cos_lut[172] = 8'hEC;
cos_lut[173] = 8'hED;
cos_lut[174] = 8'hEE;
cos_lut[175] = 8'hEF;
cos_lut[176] = 8'hF0;
cos_lut[177] = 8'hF1;
cos_lut[178] = 8'hF2;
cos_lut[179] = 8'hF3;
cos_lut[180] = 8'hF4;
cos_lut[181] = 8'hF5;
cos_lut[182] = 8'hF6;
cos_lut[183] = 8'hF7;
cos_lut[184] = 8'hF8;
cos_lut[185] = 8'hF9;
cos_lut[186] = 8'hFA;
cos_lut[187] = 8'hFB;
cos_lut[188] = 8'hFC;
cos_lut[189] = 8'hFD;
cos_lut[190] = 8'hFE;
cos_lut[191] = 8'hFF;
cos_lut[192] = 8'h00;
cos_lut[193] = 8'h01;
cos_lut[194] = 8'h02;
cos_lut[195] = 8'h03;
cos_lut[196] = 8'h04;
cos_lut[197] = 8'h05;
cos_lut[198] = 8'h06;
cos_lut[199] = 8'h07;
cos_lut[200] = 8'h08;
cos_lut[201] = 8'h09;
cos_lut[202] = 8'h0A;
cos_lut[203] = 8'h0B;
cos_lut[204] = 8'h0C;
cos_lut[205] = 8'h0D;
cos_lut[206] = 8'h0E;
cos_lut[207] = 8'h0F;
cos_lut[208] = 8'h10;
cos_lut[209] = 8'h11;
cos_lut[210] = 8'h12;
cos_lut[211] = 8'h13;
cos_lut[212] = 8'h14;
cos_lut[213] = 8'h15;
cos_lut[214] = 8'h16;
cos_lut[215] = 8'h16;
cos_lut[216] = 8'h17;
cos_lut[217] = 8'h18;
cos_lut[218] = 8'h19;
cos_lut[219] = 8'h1A;
cos_lut[220] = 8'h1B;
cos_lut[221] = 8'h1B;
cos_lut[222] = 8'h1C;
cos_lut[223] = 8'h1D;
cos_lut[224] = 8'h1E;
cos_lut[225] = 8'h1E;
cos_lut[226] = 8'h1F;
cos_lut[227] = 8'h20;
cos_lut[228] = 8'h20;
cos_lut[229] = 8'h21;
cos_lut[230] = 8'h22;
cos_lut[231] = 8'h22;
cos_lut[232] = 8'h23;
cos_lut[233] = 8'h23;
cos_lut[234] = 8'h24;
cos_lut[235] = 8'h25;
cos_lut[236] = 8'h25;
cos_lut[237] = 8'h26;
cos_lut[238] = 8'h26;
cos_lut[239] = 8'h26;
cos_lut[240] = 8'h27;
cos_lut[241] = 8'h27;
cos_lut[242] = 8'h28;
cos_lut[243] = 8'h28;
cos_lut[244] = 8'h28;
cos_lut[245] = 8'h28;
cos_lut[246] = 8'h29;
cos_lut[247] = 8'h29;
cos_lut[248] = 8'h29;
cos_lut[249] = 8'h29;
cos_lut[250] = 8'h2A;
cos_lut[251] = 8'h2A;
cos_lut[252] = 8'h2A;
cos_lut[253] = 8'h2A;
cos_lut[254] = 8'h2A;
cos_lut[255] = 8'h2A;

end

always @(posedge clock) begin
    q <= cos_lut[address];
end

endmodule
